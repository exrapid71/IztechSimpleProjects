LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
  
ENTITY REGISTER_8BIT IS PORT(
  input  : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END REGISTER_8BIT;

ARCHITECTURE BEHAVIORAL_REGISTER_8BIT OF REGISTER_8BIT IS
BEGIN
  output <= input;
END BEHAVIORAL_REGISTER_8BIT;