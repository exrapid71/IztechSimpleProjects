library ieee;
use ieee.std_logic_1164.all;

entity mux2to1 is 
port(

	
