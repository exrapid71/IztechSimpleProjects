LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU_8BIT IS PORT(
      sel :   IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      a,b :   IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      f   :  OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      unsignedOverflow : OUT STD_LOGIC;
      signedOverflow : OUT STD_LOGIC;
      carry, zero : OUT STD_LOGIC);     
END ALU_8BIT;

ARCHITECTURE ALU_8BIT_STRUCTURAL OF ALU_8BIT IS
    
    COMPONENT FA_8BIT IS PORT(
      x0, y0    :   IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      cin       :   IN STD_LOGIC;
      f         :   OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      unsignedOverflow, signedOverflow :   OUT STD_LOGIC);
    END COMPONENT;
    
    COMPONENT A_EXTENDER_8BIT IS PORT(
      s   :   IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      b   :   IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      y   :  OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
    
    COMPONENT L_EXTENDER_8BIT IS PORT(
      s   :   IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      a,b :   IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      x   :  OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
    END COMPONENT;
    
    COMPONENT SHIFTER IS PORT(
      sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
      input : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      carryOut, zer : OUT STD_LOGIC);
    END COMPONENT;
    
    COMPONENT C_EXTENDER IS PORT(
      s   :   IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      c   :   OUT STD_LOGIC);
    END COMPONENT;
    
    SIGNAL CRRY : STD_LOGIC;
    SIGNAL AR_EXT, LOG_EXT, FUL_AD : STD_LOGIC_VECTOR(7 DOWNTO 0);
    
BEGIN
    CE : C_EXTENDER PORT MAP(sel(2 DOWNTO 0), CRRY);
    LE : L_EXTENDER_8BIT PORT MAP(sel(2 DOWNTO 0), a, b, LOG_EXT);
    AE : A_EXTENDER_8BIT PORT MAP(sel(2 DOWNTO 0),b, AR_EXT);
    FA : FA_8BIT PORT MAP(LOG_EXT, AR_EXT, CRRY, FUL_AD, unsignedOverflow, signedOverflow);
    SH : SHIFTER PORT MAP(sel(4 DOWNTO 3), FUL_AD, f, carry, zero);
END ALU_8BIT_STRUCTURAL;
