LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    
ENTITY ADRESSBUS IS PORT(
   enable : IN STD_LOGIC;
   input : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
   output : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ADRESSBUS;

ARCHITECTURE BEHAVIORAL_ADRESSBUS OF ADRESSBUS IS
BEGIN
    PROCESS(enable, input)
    BEGIN
        IF(enable = '1') THEN
            output <= input;
        END IF;
    END PROCESS;
END BEHAVIORAL_ADRESSBUS;