LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
ENTITY IR_2BYTE IS PORT(
  irClk : IN STD_LOGIC;
  irLoad1 : IN STD_LOGIC;
  irLoad2 : IN STD_LOGIC;
  irReset1 : IN STD_LOGIC;
  irReset2 : IN STD_LOGIC;
  irInput : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  outputIR1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
  outputIR2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END IR_2BYTE;
ARCHITECTURE STRUCTURAL_IR_2BYTE OF IR_2BYTE IS
COMPONENT IR IS PORT(
  clk      : IN STD_LOGIC;
  irLoad   : IN STD_LOGIC;
  irReset  : IN STD_LOGIC;
  inputIR  : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  outputIR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));  
END COMPONENT;
BEGIN
  U0 : IR PORT MAP(irClk, irLoad1, irReset1, irInput, outputIR1);
  U1 : IR PORT MAP(irClk, irLoad2, irReset2, irInput, outputIR2);
END STRUCTURAL_IR_2BYTE;