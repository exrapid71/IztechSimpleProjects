library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity SHIFTER16 is port (
S:		in std_logic_vector(1 downto 0);
A:		in std_logic_vector(15 downto 0);
Y:		out std_logic_vector(15 downto 0);
carryOut:	out std_logic;
zero:		out std_logic);
end SHIFTER16;

architecture imp of SHIFTER16 is

component mux4 is port(
	S:		in std_logic_vector(1 downto 0);
	x0, x1, x2, x3: in std_logic;
	y:		out std_logic);
end component;

begin
	process(S)
	begin 
		if(S="01") then
			carryOut <= A(15);
	elsif(S="10") then
		carryOut <= A(0);
	end if;
end process;

U0:	mux4 port map(S, A(0),  '0', A(1), A(1), Y(0));
U1:	mux4 port map(S, A(1), A(0), A(2), A(2), Y(1));
U2:	mux4 port map(S, A(2), A(1), A(3), A(3), Y(2));
U3:	mux4 port map(S, A(3), A(2), A(4), A(4), Y(3));
U4:	mux4 port map(S, A(4), A(3), A(5), A(5), Y(4));
U5:	mux4 port map(S, A(5), A(4), A(6), A(6), Y(5));
U6:	mux4 port map(S, A(6), A(5), A(7), A(7), Y(6));
U7:	mux4 port map(S, A(7), A(6), A(8), A(8), Y(7));
U8:	mux4 port map(S, A(8), A(7), A(9), A(9), Y(8));
U9:	mux4 port map(S, A(9), A(8), A(10), A(10), Y(9));
U10:	mux4 port map(S, A(10), A(9), A(11), A(11), Y(10));
U11:	mux4 port map(S, A(11), A(10), A(12), A(12), Y(11));
U12:	mux4 port map(S, A(12), A(11), A(13), A(13), Y(12));
U13:	mux4 port map(S, A(13), A(12), A(14), A(14), Y(13));
U14:	mux4 port map(S, A(14), A(13), A(15), A(15), Y(14));
U15:	mux4 port map(S, A(15), A(14), '0', A(0), Y(15));

process(S)
begin 
	if(S="00")then
		if(A=0)then
			zero <= '1';
		else
			zero <= '0';
		end if;
	end if;
end process;
end imp;

