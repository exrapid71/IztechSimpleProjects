LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;

ENTITY A_EXTENDER_8BIT IS PORT(
      s   :   IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      b   :   IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      y   :  OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END A_EXTENDER_8BIT;

ARCHITECTURE A_EXTENDER_8BIT_STRUCTURAL OF A_EXTENDER_8BIT IS
    COMPONENT A_EXTENDER IS PORT(
           s   : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
           b   : IN STD_LOGIC;
           y   : OUT STD_LOGIC);
    END COMPONENT;
BEGIN
    U0 : A_EXTENDER PORT MAP(s, b(0), y(0));
    U1 : A_EXTENDER PORT MAP(s, b(1), y(1));
    U2 : A_EXTENDER PORT MAP(s, b(2), y(2));
    U3 : A_EXTENDER PORT MAP(s, b(3), y(3));
    U4 : A_EXTENDER PORT MAP(s, b(4), y(4));
    U5 : A_EXTENDER PORT MAP(s, b(5), y(5));
    U6 : A_EXTENDER PORT MAP(s, b(6), y(6));
    U7 : A_EXTENDER PORT MAP(s, b(7), y(7));
END A_EXTENDER_8BIT_STRUCTURAL;

